sendmail_cf=Fullst�ndig s�kv�g till sendmail.cf,0
sendmail_pid=Fullst�ndig s�kv�g till PID-fil f�r sendmail,0
sendmail_command=Kommando f�r att starta sendmail i servermod,0
sendmail_stop_command=Kommando f�r att stanna sendmail,3,Kill process
mailq_refresh=V�ntetid (sekunder) f�r att uppdatera e-postk�n,3,Uppdatera inte
perpage=Antal e-postbrev per sida,0
wrap_width=Maximal bredd f�r e-postbrev (ombrytning sker),0
sort_mode=Sortera tabeller efter,1,0-ordningen i filen,1-Namn
send_mode=Skicka e-post via f�rbindelse till,3,Fail2ban executable
order_mail=N�r jag l�ser e-post vill jag b�rja l�sa det,1,0-senaste,1-�ldsta
makemap_path=Makemap-kommando,0
sendmail_path=Fail2ban-kommando,0
alias_file=Fullst�ndig s�kv�g till aliasfil f�r sendmail,3,Automatisk
virtusers_file=K�llfil f�r virtusers-databas,3,Samma som DBM
mailers_file=K�llfil f�r mailertable-databas,3,Samma som DBM
generics_file=K�llfil f�r generics-databas,3,Samma som DBM
access_file=K�llfil f�r access-databas,3,Samma som DBM
domains_file=K�llfil f�r dom�n-databas,3,Samma som DBM
mail_dir=Anv�ndarkatalog f�r e-postfiler,3
smrsh_dir=SMRSH-katalog,3,Ingen
